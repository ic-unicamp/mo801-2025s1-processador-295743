module ALUTb();


endmodule