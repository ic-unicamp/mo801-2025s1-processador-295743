module ALU(
    input wire [31:0] src_a,
    input wire [31:0] src_b,
    input wire [2:0] alu_op,
    output wire [31:0] result
);


endmodule